magic
tech scmos
timestamp 1596782085
<< nwell >>
rect -9 6 21 23
<< polysilicon >>
rect 4 12 8 14
rect 4 2 8 8
rect -2 -2 8 2
rect 4 -5 8 -2
rect 4 -11 8 -9
<< ndiffusion >>
rect -6 -9 -4 -5
rect 0 -9 4 -5
rect 8 -9 12 -5
rect 16 -9 18 -5
<< pdiffusion >>
rect 0 8 4 12
rect 8 8 12 12
<< metal1 >>
rect -9 17 -4 21
rect 0 17 4 21
rect 8 17 12 21
rect 16 17 21 21
rect -4 12 0 17
rect 12 2 16 8
rect -15 -2 -6 2
rect 12 -2 27 2
rect 12 -5 16 -2
rect -4 -13 0 -9
rect -6 -17 -4 -13
rect 0 -17 4 -13
rect 8 -17 12 -13
rect 16 -17 18 -13
<< ntransistor >>
rect 4 -9 8 -5
<< ptransistor >>
rect 4 8 8 12
<< polycontact >>
rect -6 -2 -2 2
<< ndcontact >>
rect -4 -9 0 -5
rect 12 -9 16 -5
<< pdcontact >>
rect -4 8 0 12
rect 12 8 16 12
<< psubstratepcontact >>
rect -4 -17 0 -13
rect 4 -17 8 -13
rect 12 -17 16 -13
<< nsubstratencontact >>
rect -4 17 0 21
rect 4 17 8 21
rect 12 17 16 21
<< labels >>
rlabel metal1 18 19 18 19 5 vdd!
rlabel metal1 17 -15 17 -15 1 gnd!
rlabel metal1 -15 -2 -15 2 3 in
rlabel metal1 27 -2 27 2 7 out
<< end >>
