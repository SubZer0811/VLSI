magic
tech scmos
timestamp 1597235479
<< nwell >>
rect -10 16 26 30
<< polysilicon >>
rect 19 30 21 32
rect -5 23 -3 25
rect 3 23 5 25
rect -5 15 -3 19
rect 3 15 5 19
rect -5 1 -3 11
rect 3 1 5 11
rect 19 8 21 26
rect 18 4 21 8
rect 19 1 21 4
rect -5 -5 -3 -3
rect 3 -5 5 -3
rect 19 -5 21 -3
<< ndiffusion >>
rect -6 -3 -5 1
rect -3 -3 -2 1
rect 2 -3 3 1
rect 5 -3 6 1
rect 18 -3 19 1
rect 21 -3 22 1
<< pdiffusion >>
rect 18 26 19 30
rect 21 26 22 30
rect -6 19 -5 23
rect -3 19 3 23
rect 5 19 6 23
<< metal1 >>
rect -6 32 -2 36
rect 2 32 6 36
rect 10 32 18 36
rect -10 23 -6 32
rect 14 30 18 32
rect 10 19 18 23
rect -10 11 -6 15
rect 6 11 10 15
rect 14 8 18 19
rect -2 4 14 8
rect 22 15 26 26
rect 22 11 30 15
rect -2 1 2 4
rect 22 1 26 11
rect -10 -7 -6 -3
rect 6 -7 10 -3
rect 14 -7 18 -3
rect -6 -11 -2 -7
rect 2 -11 6 -7
rect 10 -11 18 -7
<< ntransistor >>
rect -5 -3 -3 1
rect 3 -3 5 1
rect 19 -3 21 1
<< ptransistor >>
rect 19 26 21 30
rect -5 19 -3 23
rect 3 19 5 23
<< polycontact >>
rect -6 11 -2 15
rect 2 11 6 15
rect 14 4 18 8
<< ndcontact >>
rect -10 -3 -6 1
rect -2 -3 2 1
rect 6 -3 10 1
rect 14 -3 18 1
rect 22 -3 26 1
<< pdcontact >>
rect 14 26 18 30
rect 22 26 26 30
rect -10 19 -6 23
rect 6 19 10 23
<< psubstratepcontact >>
rect -10 -11 -6 -7
rect -2 -11 2 -7
rect 6 -11 10 -7
<< nsubstratencontact >>
rect -10 32 -6 36
rect -2 32 2 36
rect 6 32 10 36
<< labels >>
rlabel nsubstratencontact 7 34 7 34 5 vdd
rlabel metal1 -8 13 -8 13 3 A
rlabel metal1 8 13 8 13 1 B
rlabel metal1 11 -9 11 -9 1 gnd
rlabel metal1 29 13 29 13 7 out
<< end >>
